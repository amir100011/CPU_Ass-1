-- ====================================================================
--
--	File Name:		n_bit_adder_Test.vhd
--	Description:	Test bench for 	n_bit_adder_Test 
--					
--
--	Date:			28/03/2018
--	Designer:		Amir Tsur
--
-- ====================================================================
-- Test Bench for 	n_bit_adder_Test.

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



entity 	Aritmetic_Unit_TB is
end 	Aritmetic_Unit_TB;

architecture rtl of 	Aritmetic_Unit_TB is  

component Aritmetic_Unit is generic(

  N : integer := 8
  
);

port (

  Opcode:                        in std_logic_vector(3 downto 0);--9 actions availible
  InputBusA:                     in std_logic_vector(N-1 downto 0);
  InputBusB:                     in std_logic_vector(N-1 downto 0);
  clk:                           in std_logic;
	Aritmetic_Unit_output_MUL:     out std_logic_vector(2*N-1 downto 0);
	Aritmetic_Unit_output_MAC:     out std_logic_vector(2*N-1 downto 0); 
	Aritmetic_Unit_output_MIN_MAX: out std_logic_vector(2*N-1 downto 0);
	Aritmetic_Unit_output_FA:      out std_logic_vector(2*N-1 downto 0)
		
	);-- ports declerations
end component;

signal inA_tmp,inB_tmp  : std_logic_vector(3 downto 0):=(others=>'0');
signal clk_q : std_logic:='0';
signal opcode_q : std_logic_vector(3 downto 0):=(others=>'0');
signal sum : std_logic_vector(7 downto 0):=(others=>'0');
signal mul : std_logic_vector(7 downto 0):=(others=>'0');
signal Acc : std_logic_vector(7 downto 0):=(others=>'0');
signal MIN_MAX : std_logic_vector(7 downto 0):=(others=>'0');

for tester: Aritmetic_Unit use entity work.Aritmetic_Unit;

begin
        tester : Aritmetic_Unit
        generic map (N => 4)
        port map(inputBusA=>inA_tmp, 
                 inputBusB=>inB_tmp, 
                 clk=>clk_q, 
                 Opcode=>opcode_q, 
                 Aritmetic_Unit_output_FA=>sum,
                 Aritmetic_Unit_output_MUL => mul,
                 Aritmetic_Unit_output_MAC => Acc, 
                 Aritmetic_Unit_output_MIN_MAX => MIN_MAX           
                 );
        
        testbench : process
        begin
          
          
     --TEST 0 ADD
      inA_tmp <= "0001";
      inB_tmp <= "0101";
      clk_q <= '1';
      opcode_q <= "0000";
      wait for 1 ns;
      assert(sum = "00000110") report "sum error 0" severity error;
      
      clk_q <= '0';
      wait for 1 ns;
      
      --TEST 1 MUL
      inA_tmp <= "0011";
      inB_tmp <= "0010";
      clk_q <= '1';
      opcode_q <= "0100";
      wait for 1 ns;
      assert(mul = "00000110") report "mul error 1" severity error;
      
      clk_q <= '0';
      wait for 1 ns;
      

      --TEST 2 SUB
      inA_tmp <= "0111";
      inB_tmp <= "0010";
      clk_q <= '1';
      opcode_q <= "0001";
      wait for 1 ns;
      assert(sum = "00000101") report "sum error 2" severity error;
      
      clk_q <= '0';
      wait for 1 ns;
      
      
      --TEST 3 RST
      inA_tmp <= "0001";
      inB_tmp <= "0001";
      clk_q <= '1';
      opcode_q <= "0101";
      wait for 1 ns;
      clk_q <= '0';
      wait for 1 ns;
      clk_q <= '1';
      wait for 1 ns;
      assert(Acc = "00000000") report "Acc error 3" severity error;
  
      clk_q <= '0';
      wait for 1 ns;
      
      --TEST 4 MAC
      inA_tmp <= "0110";
      inB_tmp <= "0011";
      clk_q <= '1';
      opcode_q <= "0100";
      wait for 1 ns;
      clk_q <= '0';
      wait for 1 ns;
      clk_q <= '1';
      wait for 1 ns;
      assert(Acc = "000010010") report "Acc error 4" severity error;
      
      clk_q <= '0';
      wait for 1 ns;
      
      --TEST 5 MAX
      inA_tmp <= "0111";
      inB_tmp <= "0101";
      clk_q <= '1';
      opcode_q <= "0111";
      wait for 1 ns;
      assert(MIN_MAX = "00000111") report "MIN_MAX error 5" severity error;
      
      clk_q <= '0';
      wait for 1 ns;
      
      --TEST 6 MIN
      inA_tmp <= "0010";
      inB_tmp <= "0011";
      clk_q <= '1';
      opcode_q <= "0011";
      wait for 1 ns;
      assert(MIN_MAX = "00000010") report "MIN_MAX error 6" severity error;
      
      
   end process testbench;
    
end rtl;






